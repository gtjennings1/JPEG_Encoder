module jpeg_enc_dct (
  input           clk,
  input           reset_n,
  input           dct_en,
  input  [7:0]    data_in[63:0],
  
  );
  
endmodule  